module singleadd (result, clk, set, clear);

//Output port
output result;

//Input ports
input clk, set, clear;

//Wires and Registers
wire addend, augand

