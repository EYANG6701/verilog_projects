module alu_tb;

	//Inputs are registers
	reg [15:0] a, b;
	reg [4:0] alu_code;

	//Outputs are wires
	wire [15:0] c;
	wire overflow;

	//Instantiate DUT
	alu_module DUT (
		.a(a),
		.b(b),
		.alu_code(alu_code),
		.c(c),
		.overflow(overflow)
	);

	//Testbench
	initial begin
		$display(" time |         a                 b     alu_code|         c    overflow ");
		$monitor(" %4t | %b %b %b | %b %b ", $time, a, b, alu_code, c, overflow);

		//Test cases
		//Arithmetic
		//Signed addition
		a = 16'b0000000000000000; b = 16'b0000000000000001; alu_code = 5'b00000; #15
		a = 16'b0111111100000000; b = 16'b0000001100000000; alu_code = 5'b00000; #15
	
		//Unsigned addition
		a = 16'b0000000000000000; b = 16'b0000000000000001; alu_code = 5'b00001; #15
		a = 16'b0111111100000000; b = 16'b0000001100000000; alu_code = 5'b00000; #15
	
		//Signed subtraction
		a = 16'b0000000000000000; b = 16'b0000000000000001; alu_code = 5'b00010; #15
		a = 16'b0111111100000000; b = 16'b0000001100000000; alu_code = 5'b00010; #15

		//Unisgned subtraction
		a = 16'b0000000000000000; b = 16'b0000000000000001; alu_code = 5'b00011; #15
		a = 16'b0111111100000000; b = 16'b0000001100000000; alu_code = 5'b00011; #15

		//Increment
		a = 16'b0000000000000000; b = 16'b0000000000000001; alu_code = 5'b00100; #15
		a = 16'b0111111111111111; b = 16'b0000001100000000; alu_code = 5'b00100; #15

		//Decrement
		a = 16'b0000000000000000; b = 16'b0000000000000001; alu_code = 5'b00101; #15
		a = 16'b0111111100000000; b = 16'b0000001100000000; alu_code = 5'b00101; #15

		
		//Logic
		a = 16'b1111111111111111; b = 16'b1111111111111111; alu_code = 5'b01000; #15
		a = 16'b0000000000000000; b = 16'b0000000000000000; alu_code = 5'b01000; #15
		a = 16'b1111111100000000; b = 16'b0000000011111111; alu_code = 5'b01001; #15
		a = 16'b1111111100000000; b = 16'b1111111100000000; alu_code = 5'b01000; #15
		a = 16'b1010101010101010; b = 16'b1010101010101010; alu_code = 5'b01010; #15
		a = 16'b1010101010101010; b = 16'b0000000000000000; alu_code = 5'b01100; #15

		//Shift Operation
		a = 16'b0100100100100100; b = 16'b0000000000000001; alu_code = 5'b10000; #15
		a = 16'b0100100100100100; b = 16'b0000000000000001; alu_code = 5'b10001; #15
		a = 16'b0100100100100100; b = 16'b0000000000000001; alu_code = 5'b10010; #15
		a = 16'b0100100100100100; b = 16'b0000000000000001; alu_code = 5'b10011; #15

		//Set_condition
		a = 16'b0000000000000001; b = 16'b0000000000000001; alu_code = 5'b11000; #15
		a = 16'b0000000000000000; b = 16'b0000000000000001; alu_code = 5'b11000; #15
		a = 16'b0000000000000001; b = 16'b0000000000000000; alu_code = 5'b11000; #15
		a = 16'b0000000000000001; b = 16'b0000000000000001; alu_code = 5'b11001; #15
		a = 16'b0000000000000000; b = 16'b0000000000000001; alu_code = 5'b11001; #15
		a = 16'b0000000000000001; b = 16'b0000000000000000; alu_code = 5'b11001; #15
		a = 16'b0000000000000001; b = 16'b0000000000000001; alu_code = 5'b11010; #15
		a = 16'b0000000000000000; b = 16'b0000000000000001; alu_code = 5'b11010; #15
		a = 16'b0000000000000001; b = 16'b0000000000000000; alu_code = 5'b11010; #15
		a = 16'b0000000000000001; b = 16'b0000000000000001; alu_code = 5'b11011; #15
		a = 16'b0000000000000000; b = 16'b0000000000000001; alu_code = 5'b11011; #15
		a = 16'b0000000000000001; b = 16'b0000000000000000; alu_code = 5'b11011; #15
		a = 16'b0000000000000001; b = 16'b0000000000000001; alu_code = 5'b11100; #15
		a = 16'b0000000000000000; b = 16'b0000000000000001; alu_code = 5'b11100; #15
		a = 16'b0000000000000001; b = 16'b0000000000000000; alu_code = 5'b11100; #15
		a = 16'b0000000000000001; b = 16'b0000000000000001; alu_code = 5'b11101; #15
		a = 16'b0000000000000000; b = 16'b0000000000000001; alu_code = 5'b11101; #15
		a = 16'b0000000000000001; b = 16'b0000000000000000; alu_code = 5'b11101; #15
		$finish;
	end
endmodule

	