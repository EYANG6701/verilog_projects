module csa (sum, cout, a, b, c);

    //Output ports
    output sum, cout;

    //Input ports
    input a, b, c;

    //Structural
    