module dflipflop (q, q_bar, d, clk);

    //output 
    output q, q_bar;

    //input 
    input d, clk;

    