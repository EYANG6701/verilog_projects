module alu_tb();

